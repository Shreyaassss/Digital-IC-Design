*** SPICE deck for cell FiveStageRingOsc{sch} from library Demo
*** Created on Thu Sep 05, 2024 12:41:44
*** Last revised on Thu Sep 05, 2024 14:54:58
*** Written on Thu Sep 05, 2024 17:28:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.01FF

*** SUBCIRCUIT Demo__inverter FROM CELL inverter{sch}
.SUBCKT Demo__inverter gnd INP OUT vdd
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.044U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.088U

* Spice Code nodes in cell cell 'inverter{sch}'
.include "D:\DIC\22nm_HP.pm"
.ENDS Demo__inverter

*** TOP LEVEL CELL: FiveStageRingOsc{sch}
Xinverter@0 gnd net@0 net@9 vdd Demo__inverter
Xinverter@1 gnd net@9 net@19 vdd Demo__inverter
Xinverter@2 gnd net@19 net@27 vdd Demo__inverter
Xinverter@3 gnd net@27 in1 vdd Demo__inverter
Xinverter@4 gnd in1 net@0 vdd Demo__inverter

* Spice Code nodes in cell cell 'FiveStageRingOsc{sch}'
.include "D:\DIC\22nm_HP.pm"
v1 vdd gnd DC 0.8
.ic v(in1)=0.8
.tran 0 10n 0 0.1p
.meas t1 find time when v(in1)=0.4 cross=8
.meas t2 find time when v(in1)=0.4 cross=10
.meas f param 1/(t2-t1)
.END
