*** SPICE deck for cell inverter{sch} from library Demo
*** Created on Sun Aug 18, 2024 09:29:17
*** Last revised on Mon Oct 14, 2024 21:45:27
*** Written on Mon Oct 14, 2024 21:45:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.01FF

*** TOP LEVEL CELL: inverter{sch}
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.044U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.088U

* Spice Code nodes in cell cell 'inverter{sch}'
.include "D:\DIC\22nm_HP.pm"
v1 vdd gnd DC 0.8
v2 INP gnd pwl(0 0 100p 0.8 1n 0.8 1.1n 0 2n 0)
.meas tran TPLH
.tran 2.1n
.END
.END
