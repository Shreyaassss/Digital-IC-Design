*** SPICE deck for cell Test_FA_2x{sch} from library Demo
*** Created on Thu Oct 24, 2024 16:38:56
*** Last revised on Thu Oct 24, 2024 17:53:20
*** Written on Thu Oct 24, 2024 21:30:14 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Demo__FA_2x FROM CELL FA_2x{sch}
.SUBCKT Demo__FA_2x A B C_in gnd vdd _C_out _S
Mnmos@0 _C_out C_in net@20 gnd nmos L=0.022U W=0.088U
Mnmos@1 _C_out C_in net@20 gnd nmos L=0.022U W=0.088U
Mnmos@2 net@20 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@3 net@20 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@4 net@20 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@5 net@20 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@6 _C_out A net@65 gnd nmos L=0.022U W=0.088U
Mnmos@7 net@65 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@8 _S _C_out net@92 gnd nmos L=0.022U W=0.088U
Mnmos@9 _S _C_out net@92 gnd nmos L=0.022U W=0.088U
Mnmos@10 net@92 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@11 net@92 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@12 net@92 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@13 net@92 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@14 net@92 C_in gnd gnd nmos L=0.022U W=0.088U
Mnmos@15 net@92 C_in gnd gnd nmos L=0.022U W=0.088U
Mnmos@16 net@215 B gnd gnd nmos L=0.022U W=0.066U
Mnmos@17 net@215 B gnd gnd nmos L=0.022U W=0.066U
Mnmos@18 net@227 A net@215 gnd nmos L=0.022U W=0.066U
Mnmos@19 net@227 A net@215 gnd nmos L=0.022U W=0.066U
Mnmos@20 _S C_in net@227 gnd nmos L=0.022U W=0.066U
Mnmos@21 _S C_in net@227 gnd nmos L=0.022U W=0.066U
Mpmos@0 net@0 C_in _C_out vdd pmos L=0.022U W=0.176U
Mpmos@1 net@0 C_in _C_out vdd pmos L=0.022U W=0.176U
Mpmos@2 vdd A net@0 vdd pmos L=0.022U W=0.176U
Mpmos@3 vdd A net@0 vdd pmos L=0.022U W=0.176U
Mpmos@4 vdd B net@0 vdd pmos L=0.022U W=0.176U
Mpmos@5 vdd B net@0 vdd pmos L=0.022U W=0.176U
Mpmos@6 net@55 A _C_out vdd pmos L=0.022U W=0.176U
Mpmos@7 vdd B net@55 vdd pmos L=0.022U W=0.176U
Mpmos@8 net@148 _C_out _S vdd pmos L=0.022U W=0.176U
Mpmos@9 net@148 _C_out _S vdd pmos L=0.022U W=0.176U
Mpmos@10 vdd A net@148 vdd pmos L=0.022U W=0.176U
Mpmos@11 vdd A net@148 vdd pmos L=0.022U W=0.176U
Mpmos@12 vdd B net@148 vdd pmos L=0.022U W=0.176U
Mpmos@13 vdd B net@148 vdd pmos L=0.022U W=0.176U
Mpmos@14 vdd C_in net@148 vdd pmos L=0.022U W=0.176U
Mpmos@15 vdd C_in net@148 vdd pmos L=0.022U W=0.176U
Mpmos@16 net@257 C_in _S vdd pmos L=0.022U W=0.132U
Mpmos@17 net@257 C_in _S vdd pmos L=0.022U W=0.132U
Mpmos@18 net@274 A net@257 vdd pmos L=0.022U W=0.132U
Mpmos@19 net@274 A net@257 vdd pmos L=0.022U W=0.132U
Mpmos@20 vdd B net@274 vdd pmos L=0.022U W=0.132U
Mpmos@21 vdd B net@274 vdd pmos L=0.022U W=0.132U

* Spice Code nodes in cell cell 'FA_2x{sch}'
.include "D:\DIC\22nm_HP.pm"	
.ENDS Demo__FA_2x

* cell 'inverter{sch}' is described in this file:
.include D:\DIC\inverter_RC.spi

*** TOP LEVEL CELL: Test_FA_2x{sch}
XFA_2x@2 A1 B1 C_in1 gnd vdd _C_out _S Demo__FA_2x
Xinverter@0 gnd net@75 A1 vdd Demo__inverter
Xinverter@1 gnd A net@75 vdd Demo__inverter
Xinverter@2 gnd net@86 B1 vdd Demo__inverter
Xinverter@3 gnd B net@86 vdd Demo__inverter
Xinverter@4 gnd net@91 C_in1 vdd Demo__inverter
Xinverter@5 gnd C_in net@91 vdd Demo__inverter

* Spice Code nodes in cell cell 'Test_FA_2x{sch}'
.include "D:\DIC\22nm_HP.pm"
.params vdd = 0.8
v1 vdd gnd DC {vdd}
v2 C_in gnd PWL(0 {vdd} 400p {vdd} 500p 0 0.9n 0 1n {vdd} 2.5n {vdd} )
v3 B gnd PWL(0 0 2.5n 0 )
v4 A gnd PWL(0 {vdd} 1.4n {vdd} 1.5n 0 1.9n 0 2n {vdd} 2.5n {vdd})
.meas tran tCoff
+trig v(C_in1) val={vdd/2} cross=1
+targ v(_S) val={vdd/2} cross=1
.meas tran tCon
+trig v(C_in1) val={vdd/2} cross=2
+targ v(_S) val={vdd/2} cross=2
.meas tran tAoff
+trig v(A1) val={vdd/2} cross=1
+targ v(_S) val={vdd/2} cross=3
.meas tran tAon
+trig v(A1) val={vdd/2} cross=2
+targ v(_S) val={vdd/2} cross=4
.trans 0 2.5n	
.END
