*** SPICE deck for cell Test__NAND2_2x{sch} from library Demo
*** Created on Thu Sep 26, 2024 12:55:30
*** Last revised on Thu Sep 26, 2024 15:46:07
*** Written on Thu Sep 26, 2024 15:46:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.01FF

* cell 'NAND2_2x{sch}' is described in this file:
.include D:\DIC\RC_extracted_NAND2_2x.spi

*** SUBCIRCUIT Demo__inverter FROM CELL inverter{sch}
.SUBCKT Demo__inverter gnd INP OUT vdd
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.044U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.088U

* Spice Code nodes in cell cell 'inverter{sch}'
.include "D:\DIC\22nm_HP.pm"
.ENDS Demo__inverter

*** TOP LEVEL CELL: Test__NAND2_2x{sch}
XNAND2_2x@0 A_in B_in gnd vdd Y Demo__NAND2_2x
Xinverter@0 gnd A net@8 vdd Demo__inverter
Xinverter@1 gnd net@8 A_in vdd Demo__inverter
Xinverter@2 gnd B net@15 vdd Demo__inverter
Xinverter@3 gnd net@15 B_in vdd Demo__inverter

* Spice Code nodes in cell cell 'Test__NAND2_2x{sch}'
.include "D:\DIC\22nm_HP.pm"
.params vdd = 0.8
v1 vdd gnd DC {vdd}
v2 A gnd PWL(0 0 400p 0 500p {vdd} 900p {vdd} 1n 0 1.4n 0 1.5n {vdd} 1.9n {vdd} 2n 0)
v3 B gnd PWL(0 0 900p 0 1n {vdd} 1.9n {vdd} 2n 0)
.meas tran delay_a_to_y
+trig v(a_in) val={vdd/2} cross=3
+targ v(y) val={vdd/2} cross=1
.trans 0 2n	
.END
