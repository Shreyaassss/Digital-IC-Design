*** SPICE deck for cell Test__NAND2_2x{sch} from library Demo
*** Created on Thu Sep 26, 2024 12:55:30
*** Last revised on Thu Sep 26, 2024 17:42:45
*** Written on Thu Sep 26, 2024 17:43:03 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.01FF

*** SUBCIRCUIT Demo__NAND2_2x FROM CELL NAND2_2x{sch}
.SUBCKT Demo__NAND2_2x A B gnd vdd Y
Mnmos@0 Y A net@65 gnd nmos L=0.022U W=0.176U
Mnmos@1 net@65 B gnd gnd nmos L=0.022U W=0.176U
Mpmos@0 vdd A Y vdd pmos L=0.022U W=0.176U
Mpmos@2 vdd B Y vdd pmos L=0.022U W=0.176U
.ENDS Demo__NAND2_2x

*** SUBCIRCUIT Demo__inverter FROM CELL inverter{sch}
.SUBCKT Demo__inverter gnd INP OUT vdd
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.044U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.088U

* Spice Code nodes in cell cell 'inverter{sch}'
.include "D:\DIC\22nm_HP.pm"
.ENDS Demo__inverter

*** TOP LEVEL CELL: Test__NAND2_2x{sch}
XNAND2_2x@0 A_in B_in gnd vdd Y Demo__NAND2_2x
XNAND2_2x@1 Y net@23 gnd vdd net@22 Demo__NAND2_2x
Xinverter@0 gnd A net@8 vdd Demo__inverter
Xinverter@1 gnd net@8 A_in vdd Demo__inverter
Xinverter@2 gnd B net@15 vdd Demo__inverter
Xinverter@3 gnd net@15 B_in vdd Demo__inverter

* Spice Code nodes in cell cell 'Test__NAND2_2x{sch}'
.include "D:\DIC\22nm_HP.pm"
.params vdd = 0.8
v1 vdd gnd DC {vdd}
v2 A gnd PWL(0 0 400p 0 500p {vdd} 900p {vdd} 1n 0 1.4n 0 1.5n {vdd} 1.9n {vdd} 2n 0)
v3 B gnd PWL(0 0 900p 0 1n {vdd} 1.9n {vdd})
.meas tran tPHL
+trig v(a_in) val={vdd/2} cross=3
+targ v(y) val={vdd/2} cross=1
.meas tran tPLH
+trig v(a_in) val={vdd/2} cross=4
+targ v(y) val={vdd/2} cross=2
.trans 0 2.4n
.END
