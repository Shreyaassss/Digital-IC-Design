*** SPICE deck for cell Text__FA_Carry_3x{sch} from library Demo
*** Created on Thu Oct 17, 2024 14:33:39
*** Last revised on Mon Oct 21, 2024 00:33:46
*** Written on Thu Oct 24, 2024 17:13:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Demo__FA_3x_Carry FROM CELL FA_3x_Carry{sch}
.SUBCKT Demo__FA_3x_Carry A B C_in gnd vdd _C_out
Mnmos@0 _C_out C_in net@33 gnd nmos L=0.4U W=1.6U
Mnmos@1 _C_out C_in net@33 gnd nmos L=0.4U W=1.6U
Mnmos@2 _C_out C_in net@33 gnd nmos L=0.4U W=1.6U
Mnmos@3 net@33 A gnd gnd nmos L=0.4U W=1.6U
Mnmos@4 net@33 A gnd gnd nmos L=0.4U W=1.6U
Mnmos@5 net@33 A gnd gnd nmos L=0.4U W=1.6U
Mnmos@6 net@33 B gnd gnd nmos L=0.4U W=1.6U
Mnmos@7 net@33 B gnd gnd nmos L=0.4U W=1.6U
Mnmos@8 net@33 B gnd gnd nmos L=0.4U W=1.6U
Mnmos@9 _C_out A net@18 gnd nmos L=0.4U W=1.6U
Mnmos@10 net@18 B gnd gnd nmos L=0.4U W=1.6U
Mpmos@0 net@0 C_in _C_out vdd pmos L=0.4U W=3.2U
Mpmos@1 net@0 C_in _C_out vdd pmos L=0.4U W=3.2U
Mpmos@2 net@0 C_in _C_out vdd pmos L=0.4U W=3.2U
Mpmos@3 vdd A net@0 vdd pmos L=0.4U W=3.2U
Mpmos@4 vdd A net@0 vdd pmos L=0.4U W=3.2U
Mpmos@5 vdd A net@0 vdd pmos L=0.4U W=3.2U
Mpmos@6 vdd B net@0 vdd pmos L=0.4U W=3.2U
Mpmos@7 vdd B net@0 vdd pmos L=0.4U W=3.2U
Mpmos@8 vdd B net@0 vdd pmos L=0.4U W=3.2U
Mpmos@9 net@17 A _C_out vdd pmos L=0.4U W=3.2U
Mpmos@10 vdd B net@17 vdd pmos L=0.4U W=3.2U

* Spice Code nodes in cell cell 'FA_3x_Carry{sch}'
.include "D:\DIC\22nm_HP.pm"	
.ENDS Demo__FA_3x_Carry

* cell 'inverter{sch}' is described in this file:
.include D:\DIC\inverter_RC.spi

*** TOP LEVEL CELL: Text__FA_Carry_3x{sch}
XFA_3x_Ca@0 A1 B1 C_in1 gnd vdd _C_out Demo__FA_3x_Carry
Xinverter@0 gnd A net@0 vdd Demo__inverter
Xinverter@1 gnd net@0 A1 vdd Demo__inverter
Xinverter@2 gnd B net@5 vdd Demo__inverter
Xinverter@3 gnd net@5 B1 vdd Demo__inverter
Xinverter@4 gnd C_in net@8 vdd Demo__inverter
Xinverter@5 gnd net@8 C_in1 vdd Demo__inverter
Xinverter@6 gnd _C_out net@19 vdd Demo__inverter

* Spice Code nodes in cell cell 'Text__FA_Carry_3x{sch}'
.include "D:\DIC\22nm_HP.pm"
.params vdd = 0.8
v1 vdd gnd DC {vdd}
v2 C_in gnd PWL(0 {vdd} 400p {vdd} 500p 0 0.9n 0 1n {vdd} 2.5n {vdd} )
v3 B gnd PWL(0 0 2.5n 0 )
v4 A gnd PWL(0 {vdd} 1.4n {vdd} 1.5n 0 1.9n 0 2n {vdd} 2.5n {vdd})
.meas tran tCoff
+trig v(C_in1) val={vdd/2} cross=1
+targ v(_C_out) val={vdd/2} cross=1
.meas tran tCon
+trig v(C_in1) val={vdd/2} cross=2
+targ v(_C_out) val={vdd/2} cross=2
.meas tran tAoff
+trig v(A1) val={vdd/2} cross=1
+targ v(_C_out) val={vdd/2} cross=3
.meas tran tAon
+trig v(A1) val={vdd/2} cross=2
+targ v(_C_out) val={vdd/2} cross=4
.trans 0 2.5n	
.END
